library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TEST_PLAYER_ROUND_INPUT is
    Port (  
    
        
            
            -- stdlogic outputs        
            CA    : out STD_LOGIC;     
            CB    : out STD_LOGIC;     
            CC    : out STD_LOGIC;     
            CD    : out STD_LOGIC;     
            CE    : out STD_LOGIC;     
            CF    : out STD_LOGIC;     
            CG    : out STD_LOGIC;     
            DP    : out STD_LOGIC;     
            AN1      : out STD_LOGIC;  
            AN2      : out STD_LOGIC;  
            AN3      : out STD_LOGIC;  
            AN4      : out STD_LOGIC   
    
                 );
end TEST_PLAYER_ROUND_INPUT;

architecture Behavioral of TEST_PLAYER_ROUND_INPUT is

begin


end Behavioral;
